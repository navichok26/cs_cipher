package p_table_pkg;

  // P-table lookup as a pure function (avoids array init issues in some iverilog builds).
  function automatic logic [7:0] p_lookup(input logic [7:0] din);
    case (din)
      8'h00: p_lookup = 8'h29;
      8'h01: p_lookup = 8'h0D;
      8'h02: p_lookup = 8'h61;
      8'h03: p_lookup = 8'h40;
      8'h04: p_lookup = 8'h9C;
      8'h05: p_lookup = 8'hEB;
      8'h06: p_lookup = 8'h9E;
      8'h07: p_lookup = 8'h8F;
      8'h08: p_lookup = 8'h1F;
      8'h09: p_lookup = 8'h85;
      8'h0A: p_lookup = 8'h5F;
      8'h0B: p_lookup = 8'h58;
      8'h0C: p_lookup = 8'h5B;
      8'h0D: p_lookup = 8'h01;
      8'h0E: p_lookup = 8'h39;
      8'h0F: p_lookup = 8'h86;
      8'h10: p_lookup = 8'h97;
      8'h11: p_lookup = 8'h2E;
      8'h12: p_lookup = 8'hD7;
      8'h13: p_lookup = 8'hD6;
      8'h14: p_lookup = 8'h35;
      8'h15: p_lookup = 8'hAE;
      8'h16: p_lookup = 8'h17;
      8'h17: p_lookup = 8'h16;
      8'h18: p_lookup = 8'h21;
      8'h19: p_lookup = 8'hB6;
      8'h1A: p_lookup = 8'h69;
      8'h1B: p_lookup = 8'h4E;
      8'h1C: p_lookup = 8'hA5;
      8'h1D: p_lookup = 8'h72;
      8'h1E: p_lookup = 8'h87;
      8'h1F: p_lookup = 8'h08;
      8'h20: p_lookup = 8'h3C;
      8'h21: p_lookup = 8'h18;
      8'h22: p_lookup = 8'hE6;
      8'h23: p_lookup = 8'hE7;
      8'h24: p_lookup = 8'hFA;
      8'h25: p_lookup = 8'hAD;
      8'h26: p_lookup = 8'hB8;
      8'h27: p_lookup = 8'h89;
      8'h28: p_lookup = 8'hB7;
      8'h29: p_lookup = 8'h00;
      8'h2A: p_lookup = 8'hF7;
      8'h2B: p_lookup = 8'h6F;
      8'h2C: p_lookup = 8'h73;
      8'h2D: p_lookup = 8'h84;
      8'h2E: p_lookup = 8'h11;
      8'h2F: p_lookup = 8'h63;
      8'h30: p_lookup = 8'h3F;
      8'h31: p_lookup = 8'h96;
      8'h32: p_lookup = 8'h7F;
      8'h33: p_lookup = 8'h6E;
      8'h34: p_lookup = 8'hBF;
      8'h35: p_lookup = 8'h14;
      8'h36: p_lookup = 8'h9D;
      8'h37: p_lookup = 8'hAC;
      8'h38: p_lookup = 8'hA4;
      8'h39: p_lookup = 8'h0E;
      8'h3A: p_lookup = 8'h7E;
      8'h3B: p_lookup = 8'hF6;
      8'h3C: p_lookup = 8'h20;
      8'h3D: p_lookup = 8'h4A;
      8'h3E: p_lookup = 8'h62;
      8'h3F: p_lookup = 8'h30;
      8'h40: p_lookup = 8'h03;
      8'h41: p_lookup = 8'hC5;
      8'h42: p_lookup = 8'h4B;
      8'h43: p_lookup = 8'h5A;
      8'h44: p_lookup = 8'h46;
      8'h45: p_lookup = 8'hA3;
      8'h46: p_lookup = 8'h44;
      8'h47: p_lookup = 8'h65;
      8'h48: p_lookup = 8'h7D;
      8'h49: p_lookup = 8'h4D;
      8'h4A: p_lookup = 8'h3D;
      8'h4B: p_lookup = 8'h42;
      8'h4C: p_lookup = 8'h79;
      8'h4D: p_lookup = 8'h49;
      8'h4E: p_lookup = 8'h1B;
      8'h4F: p_lookup = 8'h5C;
      8'h50: p_lookup = 8'hF5;
      8'h51: p_lookup = 8'h6C;
      8'h52: p_lookup = 8'hB5;
      8'h53: p_lookup = 8'h94;
      8'h54: p_lookup = 8'h54;
      8'h55: p_lookup = 8'hFF;
      8'h56: p_lookup = 8'h56;
      8'h57: p_lookup = 8'h57;
      8'h58: p_lookup = 8'h0B;
      8'h59: p_lookup = 8'hF4;
      8'h5A: p_lookup = 8'h43;
      8'h5B: p_lookup = 8'h0C;
      8'h5C: p_lookup = 8'h4F;
      8'h5D: p_lookup = 8'h70;
      8'h5E: p_lookup = 8'h6D;
      8'h5F: p_lookup = 8'h0A;
      8'h60: p_lookup = 8'hE4;
      8'h61: p_lookup = 8'h02;
      8'h62: p_lookup = 8'h3E;
      8'h63: p_lookup = 8'h2F;
      8'h64: p_lookup = 8'hA2;
      8'h65: p_lookup = 8'h47;
      8'h66: p_lookup = 8'hE0;
      8'h67: p_lookup = 8'hC1;
      8'h68: p_lookup = 8'hD5;
      8'h69: p_lookup = 8'h1A;
      8'h6A: p_lookup = 8'h95;
      8'h6B: p_lookup = 8'hA7;
      8'h6C: p_lookup = 8'h51;
      8'h6D: p_lookup = 8'h5E;
      8'h6E: p_lookup = 8'h33;
      8'h6F: p_lookup = 8'h2B;
      8'h70: p_lookup = 8'h5D;
      8'h71: p_lookup = 8'hD4;
      8'h72: p_lookup = 8'h1D;
      8'h73: p_lookup = 8'h2C;
      8'h74: p_lookup = 8'hEE;
      8'h75: p_lookup = 8'h75;
      8'h76: p_lookup = 8'hEC;
      8'h77: p_lookup = 8'hDD;
      8'h78: p_lookup = 8'h7C;
      8'h79: p_lookup = 8'h4C;
      8'h7A: p_lookup = 8'hA6;
      8'h7B: p_lookup = 8'hB4;
      8'h7C: p_lookup = 8'h78;
      8'h7D: p_lookup = 8'h48;
      8'h7E: p_lookup = 8'h3A;
      8'h7F: p_lookup = 8'h32;
      8'h80: p_lookup = 8'h98;
      8'h81: p_lookup = 8'hAF;
      8'h82: p_lookup = 8'hC0;
      8'h83: p_lookup = 8'hE1;
      8'h84: p_lookup = 8'h2D;
      8'h85: p_lookup = 8'h09;
      8'h86: p_lookup = 8'h0F;
      8'h87: p_lookup = 8'h1E;
      8'h88: p_lookup = 8'hB9;
      8'h89: p_lookup = 8'h27;
      8'h8A: p_lookup = 8'h8A;
      8'h8B: p_lookup = 8'hE9;
      8'h8C: p_lookup = 8'hBD;
      8'h8D: p_lookup = 8'hE3;
      8'h8E: p_lookup = 8'h9F;
      8'h8F: p_lookup = 8'h07;
      8'h90: p_lookup = 8'hB1;
      8'h91: p_lookup = 8'hEA;
      8'h92: p_lookup = 8'h92;
      8'h93: p_lookup = 8'h93;
      8'h94: p_lookup = 8'h53;
      8'h95: p_lookup = 8'h6A;
      8'h96: p_lookup = 8'h31;
      8'h97: p_lookup = 8'h10;
      8'h98: p_lookup = 8'h80;
      8'h99: p_lookup = 8'hF2;
      8'h9A: p_lookup = 8'hD8;
      8'h9B: p_lookup = 8'h9B;
      8'h9C: p_lookup = 8'h04;
      8'h9D: p_lookup = 8'h36;
      8'h9E: p_lookup = 8'h06;
      8'h9F: p_lookup = 8'h8E;
      8'hA0: p_lookup = 8'hBE;
      8'hA1: p_lookup = 8'hA9;
      8'hA2: p_lookup = 8'h64;
      8'hA3: p_lookup = 8'h45;
      8'hA4: p_lookup = 8'h38;
      8'hA5: p_lookup = 8'h1C;
      8'hA6: p_lookup = 8'h7A;
      8'hA7: p_lookup = 8'h6B;
      8'hA8: p_lookup = 8'hF3;
      8'hA9: p_lookup = 8'hA1;
      8'hAA: p_lookup = 8'hF0;
      8'hAB: p_lookup = 8'hCD;
      8'hAC: p_lookup = 8'h37;
      8'hAD: p_lookup = 8'h25;
      8'hAE: p_lookup = 8'h15;
      8'hAF: p_lookup = 8'h81;
      8'hB0: p_lookup = 8'hFB;
      8'hB1: p_lookup = 8'h90;
      8'hB2: p_lookup = 8'hE8;
      8'hB3: p_lookup = 8'hD9;
      8'hB4: p_lookup = 8'h7B;
      8'hB5: p_lookup = 8'h52;
      8'hB6: p_lookup = 8'h19;
      8'hB7: p_lookup = 8'h28;
      8'hB8: p_lookup = 8'h26;
      8'hB9: p_lookup = 8'h88;
      8'hBA: p_lookup = 8'hFC;
      8'hBB: p_lookup = 8'hD1;
      8'hBC: p_lookup = 8'hE2;
      8'hBD: p_lookup = 8'h8C;
      8'hBE: p_lookup = 8'hA0;
      8'hBF: p_lookup = 8'h34;
      8'hC0: p_lookup = 8'h82;
      8'hC1: p_lookup = 8'h67;
      8'hC2: p_lookup = 8'hDA;
      8'hC3: p_lookup = 8'hCB;
      8'hC4: p_lookup = 8'hC7;
      8'hC5: p_lookup = 8'h41;
      8'hC6: p_lookup = 8'hE5;
      8'hC7: p_lookup = 8'hC4;
      8'hC8: p_lookup = 8'hC8;
      8'hC9: p_lookup = 8'hEF;
      8'hCA: p_lookup = 8'hDB;
      8'hCB: p_lookup = 8'hC3;
      8'hCC: p_lookup = 8'hCC;
      8'hCD: p_lookup = 8'hAB;
      8'hCE: p_lookup = 8'hCE;
      8'hCF: p_lookup = 8'hED;
      8'hD0: p_lookup = 8'hD0;
      8'hD1: p_lookup = 8'hBB;
      8'hD2: p_lookup = 8'hD3;
      8'hD3: p_lookup = 8'hD2;
      8'hD4: p_lookup = 8'h71;
      8'hD5: p_lookup = 8'h68;
      8'hD6: p_lookup = 8'h13;
      8'hD7: p_lookup = 8'h12;
      8'hD8: p_lookup = 8'h9A;
      8'hD9: p_lookup = 8'hB3;
      8'hDA: p_lookup = 8'hC2;
      8'hDB: p_lookup = 8'hCA;
      8'hDC: p_lookup = 8'hDE;
      8'hDD: p_lookup = 8'h77;
      8'hDE: p_lookup = 8'hDC;
      8'hDF: p_lookup = 8'hDF;
      8'hE0: p_lookup = 8'h66;
      8'hE1: p_lookup = 8'h83;
      8'hE2: p_lookup = 8'hBC;
      8'hE3: p_lookup = 8'h8D;
      8'hE4: p_lookup = 8'h60;
      8'hE5: p_lookup = 8'hC6;
      8'hE6: p_lookup = 8'h22;
      8'hE7: p_lookup = 8'h23;
      8'hE8: p_lookup = 8'hB2;
      8'hE9: p_lookup = 8'h8B;
      8'hEA: p_lookup = 8'h91;
      8'hEB: p_lookup = 8'h05;
      8'hEC: p_lookup = 8'h76;
      8'hED: p_lookup = 8'hCF;
      8'hEE: p_lookup = 8'h74;
      8'hEF: p_lookup = 8'hC9;
      8'hF0: p_lookup = 8'hAA;
      8'hF1: p_lookup = 8'hF1;
      8'hF2: p_lookup = 8'h99;
      8'hF3: p_lookup = 8'hA8;
      8'hF4: p_lookup = 8'h59;
      8'hF5: p_lookup = 8'h50;
      8'hF6: p_lookup = 8'h3B;
      8'hF7: p_lookup = 8'h2A;
      8'hF8: p_lookup = 8'hFE;
      8'hF9: p_lookup = 8'hF9;
      8'hFA: p_lookup = 8'h24;
      8'hFB: p_lookup = 8'hB0;
      8'hFC: p_lookup = 8'hBA;
      8'hFD: p_lookup = 8'hFD;
      8'hFE: p_lookup = 8'hF8;
      8'hFF: p_lookup = 8'h55;
    endcase
  endfunction

endpackage : p_table_pkg


module p_module (
  input  logic [7:0] x,
  output logic [7:0] y
);

  always @(*) begin
    case(x[7:0]) 
      8'h00: y[7:0] = 8'h29;
      8'h01: y[7:0] = 8'h0D;
      8'h02: y[7:0] = 8'h61;
      8'h03: y[7:0] = 8'h40;
      8'h04: y[7:0] = 8'h9C;
      8'h05: y[7:0] = 8'hEB;
      8'h06: y[7:0] = 8'h9E;
      8'h07: y[7:0] = 8'h8F;
      8'h08: y[7:0] = 8'h1F;
      8'h09: y[7:0] = 8'h85;
      8'h0A: y[7:0] = 8'h5F;
      8'h0B: y[7:0] = 8'h58;
      8'h0C: y[7:0] = 8'h5B;
      8'h0D: y[7:0] = 8'h01;
      8'h0E: y[7:0] = 8'h39;
      8'h0F: y[7:0] = 8'h86;
      
      8'h10: y[7:0] = 8'h97;
      8'h11: y[7:0] = 8'h2E;
      8'h12: y[7:0] = 8'hD7;
      8'h13: y[7:0] = 8'hD6;
      8'h14: y[7:0] = 8'h35;
      8'h15: y[7:0] = 8'hAE;
      8'h16: y[7:0] = 8'h17;
      8'h17: y[7:0] = 8'h16;
      8'h18: y[7:0] = 8'h21;
      8'h19: y[7:0] = 8'hB6;
      8'h1A: y[7:0] = 8'h69;
      8'h1B: y[7:0] = 8'h4E;
      8'h1C: y[7:0] = 8'hA5;
      8'h1D: y[7:0] = 8'h72;
      8'h1E: y[7:0] = 8'h87;
      8'h1F: y[7:0] = 8'h08;

      8'h20: y[7:0] = 8'h3C;
      8'h21: y[7:0] = 8'h18;
      8'h22: y[7:0] = 8'hE6;
      8'h23: y[7:0] = 8'hE7;
      8'h24: y[7:0] = 8'hFA;
      8'h25: y[7:0] = 8'hAD;
      8'h26: y[7:0] = 8'hB8;
      8'h27: y[7:0] = 8'h89;
      8'h28: y[7:0] = 8'hB7;
      8'h29: y[7:0] = 8'h00;
      8'h2A: y[7:0] = 8'hF7;
      8'h2B: y[7:0] = 8'h6F;
      8'h2C: y[7:0] = 8'h73;
      8'h2D: y[7:0] = 8'h84;
      8'h2E: y[7:0] = 8'h11;
      8'h2F: y[7:0] = 8'h63;

      8'h30: y[7:0] = 8'h3F;
      8'h31: y[7:0] = 8'h96;
      8'h32: y[7:0] = 8'h7F;
      8'h33: y[7:0] = 8'h6E;
      8'h34: y[7:0] = 8'hBF;
      8'h35: y[7:0] = 8'h14;
      8'h36: y[7:0] = 8'h9D;
      8'h37: y[7:0] = 8'hAC;
      8'h38: y[7:0] = 8'hA4;
      8'h39: y[7:0] = 8'h0E;
      8'h3A: y[7:0] = 8'h7E;
      8'h3B: y[7:0] = 8'hF6;
      8'h3C: y[7:0] = 8'h20;
      8'h3D: y[7:0] = 8'h4A;
      8'h3E: y[7:0] = 8'h62;
      8'h3F: y[7:0] = 8'h30;

      8'h40: y[7:0] = 8'h03;
      8'h41: y[7:0] = 8'hC5;
      8'h42: y[7:0] = 8'h4B;
      8'h43: y[7:0] = 8'h5A;
      8'h44: y[7:0] = 8'h46;
      8'h45: y[7:0] = 8'hA3;
      8'h46: y[7:0] = 8'h44;
      8'h47: y[7:0] = 8'h65;
      8'h48: y[7:0] = 8'h7D;
      8'h49: y[7:0] = 8'h4D;
      8'h4A: y[7:0] = 8'h3D;
      8'h4B: y[7:0] = 8'h42;
      8'h4C: y[7:0] = 8'h79;
      8'h4D: y[7:0] = 8'h49;
      8'h4E: y[7:0] = 8'h1B;
      8'h4F: y[7:0] = 8'h5C;

      8'h50: y[7:0] = 8'hF5;
      8'h51: y[7:0] = 8'h6C;
      8'h52: y[7:0] = 8'hB5;
      8'h53: y[7:0] = 8'h94;
      8'h54: y[7:0] = 8'h54;
      8'h55: y[7:0] = 8'hFF;
      8'h56: y[7:0] = 8'h56;
      8'h57: y[7:0] = 8'h57;
      8'h58: y[7:0] = 8'h0B;
      8'h59: y[7:0] = 8'hF4;
      8'h5A: y[7:0] = 8'h43;
      8'h5B: y[7:0] = 8'h0C;
      8'h5C: y[7:0] = 8'h4F;
      8'h5D: y[7:0] = 8'h70;
      8'h5E: y[7:0] = 8'h6D;
      8'h5F: y[7:0] = 8'h0A;

      8'h60: y[7:0] = 8'hE4;
      8'h61: y[7:0] = 8'h02;
      8'h62: y[7:0] = 8'h3E;
      8'h63: y[7:0] = 8'h2F;
      8'h64: y[7:0] = 8'hA2;
      8'h65: y[7:0] = 8'h47;
      8'h66: y[7:0] = 8'hE0;
      8'h67: y[7:0] = 8'hC1;
      8'h68: y[7:0] = 8'hD5;
      8'h69: y[7:0] = 8'h1A;
      8'h6A: y[7:0] = 8'h95;
      8'h6B: y[7:0] = 8'hA7;
      8'h6C: y[7:0] = 8'h51;
      8'h6D: y[7:0] = 8'h5E;
      8'h6E: y[7:0] = 8'h33;
      8'h6F: y[7:0] = 8'h2B;

      8'h70: y[7:0] = 8'h5D;
      8'h71: y[7:0] = 8'hD4;
      8'h72: y[7:0] = 8'h1D;
      8'h73: y[7:0] = 8'h2C;
      8'h74: y[7:0] = 8'hEE;
      8'h75: y[7:0] = 8'h75;
      8'h76: y[7:0] = 8'hEC;
      8'h77: y[7:0] = 8'hDD;
      8'h78: y[7:0] = 8'h7C;
      8'h79: y[7:0] = 8'h4C;
      8'h7A: y[7:0] = 8'hA6;
      8'h7B: y[7:0] = 8'hB4;
      8'h7C: y[7:0] = 8'h78;
      8'h7D: y[7:0] = 8'h48;
      8'h7E: y[7:0] = 8'h3A;
      8'h7F: y[7:0] = 8'h32;

      8'h80: y[7:0] = 8'h98;
      8'h81: y[7:0] = 8'hAF;
      8'h82: y[7:0] = 8'hC0;
      8'h83: y[7:0] = 8'hE1;
      8'h84: y[7:0] = 8'h2D;
      8'h85: y[7:0] = 8'h09;
      8'h86: y[7:0] = 8'h0F;
      8'h87: y[7:0] = 8'h1E;
      8'h88: y[7:0] = 8'hB9;
      8'h89: y[7:0] = 8'h27;
      8'h8A: y[7:0] = 8'h8A;
      8'h8B: y[7:0] = 8'hE9;
      8'h8C: y[7:0] = 8'hBD;
      8'h8D: y[7:0] = 8'hE3;
      8'h8E: y[7:0] = 8'h9F;
      8'h8F: y[7:0] = 8'h07;

      8'h90: y[7:0] = 8'hB1;
      8'h91: y[7:0] = 8'hEA;
      8'h92: y[7:0] = 8'h92;
      8'h93: y[7:0] = 8'h93;
      8'h94: y[7:0] = 8'h53;
      8'h95: y[7:0] = 8'h6A;
      8'h96: y[7:0] = 8'h31;
      8'h97: y[7:0] = 8'h10;
      8'h98: y[7:0] = 8'h80;
      8'h99: y[7:0] = 8'hF2;
      8'h9A: y[7:0] = 8'hD8;
      8'h9B: y[7:0] = 8'h9B;
      8'h9C: y[7:0] = 8'h04;
      8'h9D: y[7:0] = 8'h36;
      8'h9E: y[7:0] = 8'h06;
      8'h9F: y[7:0] = 8'h8E;

      8'hA0: y[7:0] = 8'hBE;
      8'hA1: y[7:0] = 8'hA9;
      8'hA2: y[7:0] = 8'h64;
      8'hA3: y[7:0] = 8'h45;
      8'hA4: y[7:0] = 8'h38;
      8'hA5: y[7:0] = 8'h1C;
      8'hA6: y[7:0] = 8'h7A;
      8'hA7: y[7:0] = 8'h6B;
      8'hA8: y[7:0] = 8'hF3;
      8'hA9: y[7:0] = 8'hA1;
      8'hAA: y[7:0] = 8'hF0;
      8'hAB: y[7:0] = 8'hCD;
      8'hAC: y[7:0] = 8'h37;
      8'hAD: y[7:0] = 8'h25;
      8'hAE: y[7:0] = 8'h15;
      8'hAF: y[7:0] = 8'h81;

      8'hB0: y[7:0] = 8'hFB;
      8'hB1: y[7:0] = 8'h90;
      8'hB2: y[7:0] = 8'hE8;
      8'hB3: y[7:0] = 8'hD9;
      8'hB4: y[7:0] = 8'h7B;
      8'hB5: y[7:0] = 8'h52;
      8'hB6: y[7:0] = 8'h19;
      8'hB7: y[7:0] = 8'h28;
      8'hB8: y[7:0] = 8'h26;
      8'hB9: y[7:0] = 8'h88;
      8'hBA: y[7:0] = 8'hFC;
      8'hBB: y[7:0] = 8'hD1;
      8'hBC: y[7:0] = 8'hE2;
      8'hBD: y[7:0] = 8'h8C;
      8'hBE: y[7:0] = 8'hA0;
      8'hBF: y[7:0] = 8'h34;

      8'hC0: y[7:0] = 8'h82;
      8'hC1: y[7:0] = 8'h67;
      8'hC2: y[7:0] = 8'hDA;
      8'hC3: y[7:0] = 8'hCB;
      8'hC4: y[7:0] = 8'hC7;
      8'hC5: y[7:0] = 8'h41;
      8'hC6: y[7:0] = 8'hE5;
      8'hC7: y[7:0] = 8'hC4;
      8'hC8: y[7:0] = 8'hC8;
      8'hC9: y[7:0] = 8'hEF;
      8'hCA: y[7:0] = 8'hDB;
      8'hCB: y[7:0] = 8'hC3;
      8'hCC: y[7:0] = 8'hCC;
      8'hCD: y[7:0] = 8'hAB;
      8'hCE: y[7:0] = 8'hCE;
      8'hCF: y[7:0] = 8'hED;

      8'hD0: y[7:0] = 8'hD0;
      8'hD1: y[7:0] = 8'hBB;
      8'hD2: y[7:0] = 8'hD3;
      8'hD3: y[7:0] = 8'hD2;
      8'hD4: y[7:0] = 8'h71;
      8'hD5: y[7:0] = 8'h68;
      8'hD6: y[7:0] = 8'h13;
      8'hD7: y[7:0] = 8'h12;
      8'hD8: y[7:0] = 8'h9A;
      8'hD9: y[7:0] = 8'hB3;
      8'hDA: y[7:0] = 8'hC2;
      8'hDB: y[7:0] = 8'hCA;
      8'hDC: y[7:0] = 8'hDE;
      8'hDD: y[7:0] = 8'h77;
      8'hDE: y[7:0] = 8'hDC;
      8'hDF: y[7:0] = 8'hDF;

      8'hE0: y[7:0] = 8'h66;
      8'hE1: y[7:0] = 8'h83;
      8'hE2: y[7:0] = 8'hBC;
      8'hE3: y[7:0] = 8'h8D;
      8'hE4: y[7:0] = 8'h60;
      8'hE5: y[7:0] = 8'hC6;
      8'hE6: y[7:0] = 8'h22;
      8'hE7: y[7:0] = 8'h23;
      8'hE8: y[7:0] = 8'hB2;
      8'hE9: y[7:0] = 8'h8B;
      8'hEA: y[7:0] = 8'h91;
      8'hEB: y[7:0] = 8'h05;
      8'hEC: y[7:0] = 8'h76;
      8'hED: y[7:0] = 8'hCF;
      8'hEE: y[7:0] = 8'h74;
      8'hEF: y[7:0] = 8'hC9;      

      8'hF0: y[7:0] = 8'hAA;
      8'hF1: y[7:0] = 8'hF1;
      8'hF2: y[7:0] = 8'h99;
      8'hF3: y[7:0] = 8'hA8;
      8'hF4: y[7:0] = 8'h59;
      8'hF5: y[7:0] = 8'h50;
      8'hF6: y[7:0] = 8'h3B;
      8'hF7: y[7:0] = 8'h2A;
      8'hF8: y[7:0] = 8'hFE;
      8'hF9: y[7:0] = 8'hF9;
      8'hFA: y[7:0] = 8'h24;
      8'hFB: y[7:0] = 8'hB0;
      8'hFC: y[7:0] = 8'hBA;
      8'hFD: y[7:0] = 8'hFD;
      8'hFE: y[7:0] = 8'hF8;
      8'hFF: y[7:0] = 8'h55;   
    endcase
  end

endmodule

